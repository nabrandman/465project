module xor1 (input a, input b, output y);

    xor(y, a,b);

endmodule
