module or1 (input a, input b, output y);
    //same as w/ the and this is basically just for consistencies sake
    or(y, a,b);

endmodule
